module HDU (
    input [3:0] SRC1_IN, SRC2_IN, Dest_EXE_IN, Dest_MEM_IN,
    input WB_EN_EXE, WB_EN_MEM,
    
    output hazard

);
    
endmodule